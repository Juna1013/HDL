module display_test;
