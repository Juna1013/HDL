module blink_led (
    input CLK100MHZ,
    output LED
);
